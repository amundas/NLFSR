`ifndef _build_settings_vh_
`define _build_settings_vh_

    `define SHIFTREG_WIDTH 32
    `define NUM_NLIN 1
    `define NUM_NLIN_IDX 2
    `define NUM_TESTERS 50
    `define BRANCHES_PER_LEVEL 5

    `define REF_CLK_FREQ 200e6
    `define CLK_MULT 6
    `define FAST_CLK_DIV 3.5
    `define SLOW_CLK_DIV 6

    `define UART_BAUD 2_000_000

`endif